----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    00:01:24 07/12/2025 
-- Design Name: 
-- Module Name:    full_adder_struct - Structural
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity full_adder_struct is
    Port (
        a     : in  std_logic;
        b     : in  std_logic;
        cin   : in  std_logic;
        sum   : out std_logic;
        cout  : out std_logic
    );
end full_adder_struct;

architecture Structural of full_adder_struct is

    signal s1, c1, c2 : std_logic;

    component half_adder
        Port (
            a     : in  std_logic;
            b     : in  std_logic;
            sum   : out std_logic;
            carry : out std_logic
        );
    end component;

begin
    HA1: half_adder port map(a => a,    b => b,    sum => s1, carry => c1);
    HA2: half_adder port map(a => s1,   b => cin,  sum => sum, carry => c2);
    cout <= c1 or c2;
end Structural;

